module stack (
);
    
endmodule