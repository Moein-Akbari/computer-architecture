module controller (

);
    
endmodule