module eight_queen (
);
    
endmodule