module datapath (
    // bus_in,
    // shift_to_right,
    // shift_to_left,
    // column_out
);
    // input bus_in[0:2];
    // input shift_to_left, shift_to_right;
    // output bus_out[0:2];
endmodule