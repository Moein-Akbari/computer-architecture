module eight_queen (
    start, 
    reset, 
    ready,
    out_bus);
    input start, reset;
    output ready;
    output [7:0] out_bus;
    
    controller

endmodule