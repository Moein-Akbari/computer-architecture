module stacked_controller (

);


endmodule