// module increamenter_testbench ();
//     reg enable_output,
//     reg in,
//     out,
//     carry_out
// endmodule