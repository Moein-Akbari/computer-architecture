module stack (
    clk,
    reset,
    push,
    in_data,
    pop,
    out_data,
    enable_output
); 

endmodule